///////////////////////////////////////////////
// file name  : my_interface.sv
// creat time : 2020-04-11
// author     : Gong Yingfan
// version    : v1.0
// descript   : my_interface.sv
// log        : no
///////////////////////////////////////////////

//  Interface: my_interface
//
interface my_interface
    /*  package imports  */
    #(
        // parameter_list
    )(
        // port_list
    );


    // DUT ports

    // clocking block
    
    // assert and cover property

    // other tasks and functions
    
endinterface: my_interface
