// Clock Period, default: 10ns
`ifndef PERIOD
`define PERIOD 10
`endif

// simulation timeout, default: 5s
`ifndef TIMEOUT
`define TIMEOUT 5s
`endif

// DUT parameters
